`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/07/23 22:39:37
// Design Name: 
// Module Name: data
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module data(
input clk,clr,move,store,start,
input u,d,l,r,
output reg move_able,
output [199:0] data_out
    );
    
reg       [4:0] n,n_r1,n_r2,n_r3;
reg       [3:0] m,m_r1,m_r2,m_r3;
reg       [6:0] block;
reg [9:0] R [19:0];


assign data_out = {R[19],R[18],R[17],R[16],R[15],R[14],R[13],R[12],R[11],R[10],R[9],R[8],R[7],R[6],R[5],R[4],R[3],R[2],R[1],R[0]};

always @(posedge clk)
    begin
        if (clr)begin 
        n_r1 <= 0;
        m_r1 <= 0;
        n_r2 <= 0;
        m_r2 <= 0;
        n_r3 <= 0;
        m_r3 <= 0;
        end       
        else begin
        n_r1 <= n;
        n_r2 <= n_r1;
        n_r3 <= n_r2;
        m_r1 <= m;
        m_r2 <= m_r1;
        m_r3 <= m_r2;
        end
        end
        
always @ (*)
    begin
    if (u)
        begin
            if(n>=1)begin
                if (!(R[n-1][m]))
                    move_able=1;
                else move_able=0;    
                    end
            else move_able=0;
        end
    else if (l)  
            begin
                if (m>=1)begin
                     if (!(R[n][m-1]))
                        move_able=1;
                     else move_able=0;   
                        end
                else move_able=0;         
            end          
    else if (r)  
            begin
                if (m<=8)begin
                     if (!(R[n][m+1]))
                        move_able=1;
                     else move_able=0;   
                        end
                else move_able=0;         
            end                       
    else if (d)  
            begin
                if (n<=22)begin
                     if (!(R[n+1][m]))
                        move_able=1;
                     else move_able=0;   
                        end
                else move_able=0;         
            end
         end 
         

 integer i,j;
    always @ (posedge clk or posedge clr)
    begin
        if (clr)
            begin
             R[n][m]<=1; R[0][1]<=0; R[0][2]<=0; R[0][3]<=0; R[0][4]<=0; R[0][5]<=0; R[0][6]<=0; R[0][7]<=0; R[0][8]<=0; R[0][9]<=0;
             R[1][0]<=0; R[1][1]<=0; R[1][2]<=0; R[1][3]<=0; R[1][4]<=0; R[1][5]<=0; R[1][6]<=0; R[1][7]<=0; R[1][8]<=0; R[1][9]<=0;
             R[2][0]<=0; R[2][1]<=0; R[2][2]<=0; R[2][3]<=0; R[2][4]<=0; R[2][5]<=0; R[2][6]<=0; R[2][7]<=0; R[2][8]<=0; R[2][9]<=0;
             R[3][0]<=0; R[3][1]<=0; R[3][2]<=0; R[3][3]<=0; R[3][4]<=0; R[3][5]<=0; R[3][6]<=0; R[3][7]<=0; R[3][8]<=0; R[3][9]<=0;
             R[4][0]<=0; R[4][1]<=0; R[4][2]<=0; R[4][3]<=0; R[4][4]<=0; R[4][5]<=0; R[4][6]<=0; R[4][7]<=0; R[4][8]<=0; R[4][9]<=0;
             R[5][0]<=0; R[5][1]<=0; R[5][2]<=0; R[5][3]<=0; R[5][4]<=0; R[5][5]<=0; R[5][6]<=0; R[5][7]<=0; R[5][8]<=0; R[5][9]<=0;
             R[6][0]<=0; R[6][1]<=0; R[6][2]<=0; R[6][3]<=0; R[6][4]<=0; R[6][5]<=0; R[6][6]<=0; R[6][7]<=0; R[6][8]<=0; R[6][9]<=0;           
             R[7][0]<=0; R[7][1]<=0; R[7][2]<=0; R[7][3]<=0; R[7][4]<=0; R[7][5]<=0; R[7][6]<=0; R[7][7]<=0; R[7][8]<=0; R[7][9]<=0;   
             R[8][0]<=0; R[8][1]<=0; R[8][2]<=0; R[8][3]<=0; R[8][4]<=0; R[8][5]<=0; R[8][6]<=0; R[8][7]<=0; R[8][8]<=0; R[8][9]<=0;   
             R[9][0]<=0; R[9][1]<=0; R[9][2]<=0; R[9][3]<=0; R[9][4]<=0; R[9][5]<=0; R[9][6]<=0; R[9][7]<=0; R[9][8]<=0; R[9][9]<=0;   
             R[10][0]<=0; R[10][1]<=0; R[10][2]<=0; R[10][3]<=1; R[10][4]<=1; R[10][5]<=1; R[10][6]<=1; R[10][7]<=0; R[10][8]<=0; R[10][9]<=0;   
             R[11][0]<=0; R[11][1]<=0; R[11][2]<=0; R[11][3]<=0; R[11][4]<=0; R[11][5]<=0; R[11][6]<=0; R[11][7]<=0; R[11][8]<=0; R[11][9]<=0;
             R[12][0]<=0; R[12][1]<=0; R[12][2]<=0; R[12][3]<=0; R[12][4]<=0; R[12][5]<=0; R[12][6]<=0; R[12][7]<=0; R[12][8]<=0; R[12][9]<=0;   
             R[13][0]<=0; R[13][1]<=0; R[13][2]<=0; R[13][3]<=0; R[13][4]<=0; R[13][5]<=0; R[13][6]<=0; R[13][7]<=0; R[13][8]<=0; R[13][9]<=0;
             R[14][0]<=0; R[14][1]<=0; R[14][2]<=0; R[14][3]<=0; R[14][4]<=0; R[14][5]<=0; R[14][6]<=0; R[14][7]<=0; R[14][8]<=0; R[14][9]<=0;
             R[15][0]<=0; R[15][1]<=0; R[15][2]<=0; R[15][3]<=0; R[15][4]<=0; R[15][5]<=0; R[15][6]<=0; R[15][7]<=0; R[15][8]<=0; R[15][9]<=0;
             R[16][0]<=0; R[16][1]<=0; R[16][2]<=0; R[16][3]<=0; R[16][4]<=0; R[16][5]<=0; R[16][6]<=0; R[16][7]<=0; R[16][8]<=0; R[16][9]<=0;
             R[17][0]<=0; R[17][1]<=0; R[17][2]<=0; R[17][3]<=0; R[17][4]<=0; R[17][5]<=0; R[17][6]<=0; R[17][7]<=0; R[17][8]<=0; R[17][9]<=0;
             R[18][0]<=0; R[18][1]<=0; R[18][2]<=0; R[18][3]<=0; R[18][4]<=0; R[18][5]<=0; R[18][6]<=0; R[18][7]<=0; R[18][8]<=0; R[18][9]<=0;
             R[19][0]<=0; R[19][1]<=0; R[19][2]<=0; R[19][3]<=0; R[19][4]<=0; R[19][5]<=0; R[19][6]<=0; R[19][7]<=0; R[19][8]<=0; R[19][9]<=0;              
            end                
        else if (store)
        begin
             R[n][m]<=1;
             R[n_r2][m_r2]<=0;
             R[n_r3][m_r3]<=0;
        end
         else
                R[n][m]<=R[n][m];
      end

 always @ (posedge clk or posedge clr)
    begin
        if (clr)
            n <= 0;
        else if ((move_able)&(d))
            n <= n+1;
        else if ((move_able)&(u))
            n <= n-1;
        else
            n <= n;
    end
  
  always @ (posedge clk or posedge clr)
    begin
        if (clr)
            m <= 0;
        else if  ((move_able)&(l))
             m <= m-1;
        else if  ((move_able)&(r))
             m <= m+1;
        else
            m <= m;
    end
                          
endmodule
