`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/07/23 22:39:37
// Design Name: 
// Module Name: data
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module data(
input clk,clr,move,store,start,judge,vga_control,U,D,L,R,
output reg move_able,judge_able,
output [799:0] data_b,data_q
    );
    
reg       [5:0] n,n_r1,n_r2,n_r3,n_r4;
reg       [5:0] m,m_r1,m_r2,m_r3,m_r4;
reg       [6:0] block;
reg       [19:0] R_b [39:0];
reg       [19:0] R_q [39:0];
reg test;
reg       u_r,d_r,l_r,r_r;

assign data_b = {R_b[39],R_b[38],R_b[37],R_b[36],R_b[35],R_b[34],R_b[33],R_b[32],R_b[31],R_b[30],R_b[29],R_b[28],R_b[27],R_b[26],R_b[25],R_b[24],R_b[23],R_b[22],R_b[21],R_b[20],R_b[19],R_b[18],R_b[17],R_b[16],R_b[15],R_b[14],R_b[13],R_b[12],R_b[11],R_b[10],R_b[9],R_b[8],R_b[7],R_b[6],R_b[5],R_b[4],R_b[3],R_b[2],R_b[1],R_b[0]};
assign data_q = {R_q[39],R_q[38],R_q[37],R_q[36],R_q[35],R_q[34],R_q[33],R_q[32],R_q[31],R_q[30],R_q[29],R_q[28],R_q[27],R_q[26],R_q[25],R_q[24],R_q[23],R_q[22],R_q[21],R_q[20],R_q[19],R_q[18],R_q[17],R_q[16],R_q[15],R_q[14],R_q[13],R_q[12],R_q[11],R_q[10],R_q[9],R_q[8],R_q[7],R_q[6],R_q[5],R_q[4],R_q[3],R_q[2],R_q[1],R_q[0]};

always @(posedge clk)
    begin
        if (clr)begin 
        n_r1 <= 0;
        m_r1 <= 0;
        n_r2 <= 0;
        m_r2 <= 0;
        r_r  <= 0;
        l_r  <= 0;
        u_r  <= 0;
        d_r  <= 0;
        end       
        else begin
        n_r1 <= n;
        n_r2 <= n_r1;
        m_r1 <= m;
        m_r2 <= m_r1;
        r_r  <= R;
        l_r  <= L;
        u_r  <= U;
        d_r  <= D;
        end
        end
        
always @ (*)
    begin
    move_able=0;
    if (move)begin
    if (u_r)
        begin
            if(n>0)begin
                if ((R_b[n-1][m])==0)
                    move_able=1;
                else if((R_b[n-1][m])==1)
                move_able=0;    
                    end
            else move_able=0;
        end
    else if (l_r)  
            begin
                if (m>0)begin
                     if ((R_b[n][m-1])==0)
                        move_able=1;
                     else if ((R_b[n][m-1])==1)  
                     move_able=0;   
                        end
                else move_able=0;         
            end          
    else if (r_r)  
            begin
                if (m<19)begin
                     if ((R_b[n][m+1])==0)
                        move_able=1;
                     else if ((R_b[n][m+1])==1)
                     move_able=0;   
                        end
                else move_able=0;         
            end                       
    else if (d_r)  
            begin
                if (n<39)begin
                     if ((R_b[n+1][m])==0)
                        move_able=1;
                     else if ((R_b[n+1][m])==1)
                      move_able=0;   
                        end
                else move_able=0;         
            end
         end 
       end  

    always @ (posedge clk or posedge clr)
    begin
        if (clr)
            begin
             R_b[n][m]<=1; R_b[0][1]<=0; R_b[0][2]<=0; R_b[0][3]<=1; R_b[0][4]<=0; R_b[0][5]<=0; R_b[0][6]<=0; R_b[0][7]<=1; R_b[0][8]<=1; R_b[0][9]<=1;R_b[0][10]<=1; R_b[0][11]<=0; R_b[0][12]<=0; R_b[0][13]<=0; R_b[0][14]<=0; R_b[0][15]<=0; R_b[0][16]<=0; R_b[0][17]<=0; R_b[0][18]<=0; R_b[0][19]<=0;
             R_b[1][0]<=0; R_b[1][1]<=0; R_b[1][2]<=0; R_b[1][3]<=1; R_b[1][4]<=0; R_b[1][5]<=0; R_b[1][6]<=0; R_b[1][7]<=0; R_b[1][8]<=0; R_b[1][9]<=0;R_b[1][10]<=0; R_b[1][11]<=0; R_b[1][12]<=0; R_b[1][13]<=0; R_b[1][14]<=1; R_b[1][15]<=1; R_b[1][16]<=1; R_b[1][17]<=1; R_b[1][18]<=1; R_b[1][19]<=0;
             R_b[2][0]<=0; R_b[2][1]<=0; R_b[2][2]<=0; R_b[2][3]<=1; R_b[2][4]<=1; R_b[2][5]<=0; R_b[2][6]<=0; R_b[2][7]<=0; R_b[2][8]<=0; R_b[2][9]<=0;R_b[2][10]<=0; R_b[2][11]<=0; R_b[2][12]<=0; R_b[2][13]<=0; R_b[2][14]<=0; R_b[2][15]<=0; R_b[2][16]<=0; R_b[2][17]<=0; R_b[2][18]<=1; R_b[2][19]<=0;
             R_b[3][0]<=0; R_b[3][1]<=0; R_b[3][2]<=0; R_b[3][3]<=0; R_b[3][4]<=0; R_b[3][5]<=0; R_b[3][6]<=0; R_b[3][7]<=1; R_b[3][8]<=1; R_b[3][9]<=1;R_b[3][10]<=0; R_b[3][11]<=0; R_b[3][12]<=0; R_b[3][13]<=0; R_b[3][14]<=0; R_b[3][15]<=1; R_b[3][16]<=1; R_b[3][17]<=0; R_b[3][18]<=0; R_b[3][19]<=0;
             R_b[4][0]<=1; R_b[4][1]<=0; R_b[4][2]<=0; R_b[4][3]<=0; R_b[4][4]<=0; R_b[4][5]<=0; R_b[4][6]<=0; R_b[4][7]<=0; R_b[4][8]<=0; R_b[4][9]<=1;R_b[4][10]<=0; R_b[4][11]<=0; R_b[4][12]<=0; R_b[4][13]<=0; R_b[4][14]<=0; R_b[4][15]<=0; R_b[4][16]<=0; R_b[4][17]<=0; R_b[4][18]<=0; R_b[4][19]<=0;
             R_b[5][0]<=1; R_b[5][1]<=1; R_b[5][2]<=1; R_b[5][3]<=1; R_b[5][4]<=0; R_b[5][5]<=0; R_b[5][6]<=0; R_b[5][7]<=0; R_b[5][8]<=0; R_b[5][9]<=1;R_b[5][10]<=0; R_b[5][11]<=1; R_b[5][12]<=1; R_b[5][13]<=0; R_b[5][14]<=1; R_b[5][15]<=0; R_b[5][16]<=0; R_b[5][17]<=0; R_b[5][18]<=0; R_b[5][19]<=0;
             R_b[6][0]<=1; R_b[6][1]<=0; R_b[6][2]<=0; R_b[6][3]<=0; R_b[6][4]<=0; R_b[6][5]<=0; R_b[6][6]<=0; R_b[6][7]<=0; R_b[6][8]<=0; R_b[6][9]<=1;R_b[6][10]<=0; R_b[6][11]<=0; R_b[6][12]<=0; R_b[6][13]<=0; R_b[6][14]<=1; R_b[6][15]<=0; R_b[6][16]<=0; R_b[6][17]<=1; R_b[6][18]<=1; R_b[6][19]<=0;           
             R_b[7][0]<=0; R_b[7][1]<=0; R_b[7][2]<=0; R_b[7][3]<=0; R_b[7][4]<=0; R_b[7][5]<=0; R_b[7][6]<=1; R_b[7][7]<=1; R_b[7][8]<=0; R_b[7][9]<=0;R_b[7][10]<=0; R_b[7][11]<=0; R_b[7][12]<=0; R_b[7][13]<=0; R_b[7][14]<=1; R_b[7][15]<=0; R_b[7][16]<=0; R_b[7][17]<=0; R_b[7][18]<=0; R_b[7][19]<=0;   
             R_b[8][0]<=0; R_b[8][1]<=0; R_b[8][2]<=0; R_b[8][3]<=0; R_b[8][4]<=0; R_b[8][5]<=0; R_b[8][6]<=0; R_b[8][7]<=0; R_b[8][8]<=0; R_b[8][9]<=0;R_b[8][10]<=0; R_b[8][11]<=0; R_b[8][12]<=0; R_b[8][13]<=0; R_b[8][14]<=1; R_b[8][15]<=0; R_b[8][16]<=0; R_b[8][17]<=0; R_b[8][18]<=0; R_b[8][19]<=0;   
             R_b[9][0]<=0; R_b[9][1]<=0; R_b[9][2]<=0; R_b[9][3]<=0; R_b[9][4]<=0; R_b[9][5]<=0; R_b[9][6]<=0; R_b[9][7]<=1; R_b[9][8]<=0; R_b[9][9]<=0;R_b[9][10]<=1; R_b[9][11]<=0; R_b[9][12]<=0; R_b[9][13]<=0; R_b[9][14]<=1; R_b[9][15]<=1; R_b[9][16]<=1; R_b[9][17]<=0; R_b[9][18]<=0; R_b[9][19]<=0;   
             R_b[10][0]<=0; R_b[10][1]<=1; R_b[10][2]<=1; R_b[10][3]<=1; R_b[10][4]<=1; R_b[10][5]<=0; R_b[10][6]<=0; R_b[10][7]<=1; R_b[10][8]<=0; R_b[10][9]<=0;R_b[10][10]<=1; R_b[10][11]<=0; R_b[10][12]<=0; R_b[10][13]<=0; R_b[10][14]<=0; R_b[10][15]<=0; R_b[10][16]<=0; R_b[10][17]<=0; R_b[10][18]<=0; R_b[10][19]<=1;   
             R_b[11][0]<=0; R_b[11][1]<=1; R_b[11][2]<=0; R_b[11][3]<=0; R_b[11][4]<=0; R_b[11][5]<=0; R_b[11][6]<=0; R_b[11][7]<=0; R_b[11][8]<=0; R_b[11][9]<=0;R_b[11][10]<=1; R_b[11][11]<=0; R_b[11][12]<=0; R_b[11][13]<=0; R_b[11][14]<=0; R_b[11][15]<=0; R_b[11][16]<=0; R_b[11][17]<=0; R_b[11][18]<=0; R_b[11][19]<=1;
             R_b[12][0]<=0; R_b[12][1]<=1; R_b[12][2]<=0; R_b[12][3]<=0; R_b[12][4]<=0; R_b[12][5]<=0; R_b[12][6]<=0; R_b[12][7]<=0; R_b[12][8]<=0; R_b[12][9]<=0;R_b[12][10]<=0; R_b[12][11]<=0; R_b[12][12]<=0; R_b[12][13]<=1; R_b[12][14]<=1; R_b[12][15]<=0; R_b[12][16]<=0; R_b[12][17]<=0; R_b[12][18]<=0; R_b[12][19]<=1;   
             R_b[13][0]<=0; R_b[13][1]<=0; R_b[13][2]<=0; R_b[13][3]<=0; R_b[13][4]<=1; R_b[13][5]<=1; R_b[13][6]<=1; R_b[13][7]<=1; R_b[13][8]<=1; R_b[13][9]<=0;R_b[13][10]<=0; R_b[13][11]<=0; R_b[13][12]<=0; R_b[13][13]<=0; R_b[13][14]<=0; R_b[13][15]<=0; R_b[13][16]<=0; R_b[13][17]<=0; R_b[13][18]<=0; R_b[13][19]<=1;
             R_b[14][0]<=0; R_b[14][1]<=0; R_b[14][2]<=0; R_b[14][3]<=0; R_b[14][4]<=0; R_b[14][5]<=0; R_b[14][6]<=0; R_b[14][7]<=0; R_b[14][8]<=0; R_b[14][9]<=0;R_b[14][10]<=0; R_b[14][11]<=0; R_b[14][12]<=0; R_b[14][13]<=0; R_b[14][14]<=0; R_b[14][15]<=0; R_b[14][16]<=1; R_b[14][17]<=1; R_b[14][18]<=1; R_b[14][19]<=1;
             R_b[15][0]<=0; R_b[15][1]<=0; R_b[15][2]<=0; R_b[15][3]<=0; R_b[15][4]<=0; R_b[15][5]<=0; R_b[15][6]<=0; R_b[15][7]<=0; R_b[15][8]<=0; R_b[15][9]<=0;R_b[15][10]<=0; R_b[15][11]<=1; R_b[15][12]<=1; R_b[15][13]<=1; R_b[15][14]<=1; R_b[15][15]<=0; R_b[15][16]<=0; R_b[15][17]<=0; R_b[15][18]<=0; R_b[15][19]<=0;
             R_b[16][0]<=0; R_b[16][1]<=0; R_b[16][2]<=0; R_b[16][3]<=0; R_b[16][4]<=1; R_b[16][5]<=1; R_b[16][6]<=0; R_b[16][7]<=0; R_b[16][8]<=0; R_b[16][9]<=0;R_b[16][10]<=0; R_b[16][11]<=0; R_b[16][12]<=0; R_b[16][13]<=0; R_b[16][14]<=0; R_b[16][15]<=0; R_b[16][16]<=0; R_b[16][17]<=0; R_b[16][18]<=0; R_b[16][19]<=0;
             R_b[17][0]<=0; R_b[17][1]<=0; R_b[17][2]<=1; R_b[17][3]<=0; R_b[17][4]<=0; R_b[17][5]<=0; R_b[17][6]<=0; R_b[17][7]<=0; R_b[17][8]<=0; R_b[17][9]<=0;R_b[17][10]<=0; R_b[17][11]<=0; R_b[17][12]<=0; R_b[17][13]<=0; R_b[17][14]<=0; R_b[17][15]<=0; R_b[17][16]<=0; R_b[17][17]<=0; R_b[17][18]<=0; R_b[17][19]<=0;
             R_b[18][0]<=1; R_b[18][1]<=0; R_b[18][2]<=1; R_b[18][3]<=0; R_b[18][4]<=0; R_b[18][5]<=0; R_b[18][6]<=1; R_b[18][7]<=1; R_b[18][8]<=1; R_b[18][9]<=0;R_b[18][10]<=0; R_b[18][11]<=0; R_b[18][12]<=0; R_b[18][13]<=0; R_b[18][14]<=1; R_b[18][15]<=1; R_b[18][16]<=1; R_b[18][17]<=1; R_b[18][18]<=0; R_b[18][19]<=0;
             R_b[19][0]<=1; R_b[19][1]<=0; R_b[19][2]<=1; R_b[19][3]<=0; R_b[19][4]<=0; R_b[19][5]<=0; R_b[19][6]<=0; R_b[19][7]<=0; R_b[19][8]<=1; R_b[19][9]<=0;R_b[19][10]<=0; R_b[19][11]<=1; R_b[19][12]<=0; R_b[19][13]<=0; R_b[19][14]<=0; R_b[19][15]<=0; R_b[19][16]<=0; R_b[19][17]<=0; R_b[19][18]<=0; R_b[19][19]<=0;
             R_b[20][0]<=0; R_b[20][1]<=0; R_b[20][2]<=1; R_b[20][3]<=0; R_b[20][4]<=0; R_b[20][5]<=0; R_b[20][6]<=0; R_b[20][7]<=0; R_b[20][8]<=1; R_b[20][9]<=0;R_b[20][10]<=0; R_b[20][11]<=1; R_b[20][12]<=0; R_b[20][13]<=0; R_b[20][14]<=0; R_b[20][15]<=0; R_b[20][16]<=0; R_b[20][17]<=0; R_b[20][18]<=0; R_b[20][19]<=0;   
             R_b[21][0]<=0; R_b[21][1]<=0; R_b[21][2]<=1; R_b[21][3]<=0; R_b[21][4]<=0; R_b[21][5]<=0; R_b[21][6]<=0; R_b[21][7]<=0; R_b[21][8]<=0; R_b[21][9]<=0;R_b[21][10]<=0; R_b[21][11]<=0; R_b[21][12]<=0; R_b[21][13]<=0; R_b[21][14]<=0; R_b[21][15]<=0; R_b[21][16]<=0; R_b[21][17]<=0; R_b[21][18]<=1; R_b[21][19]<=0;
             R_b[22][0]<=0; R_b[22][1]<=0; R_b[22][2]<=0; R_b[22][3]<=0; R_b[22][4]<=0; R_b[22][5]<=0; R_b[22][6]<=0; R_b[22][7]<=0; R_b[22][8]<=0; R_b[22][9]<=0;R_b[22][10]<=0; R_b[22][11]<=0; R_b[22][12]<=0; R_b[22][13]<=0; R_b[22][14]<=0; R_b[22][15]<=0; R_b[22][16]<=0; R_b[22][17]<=0; R_b[22][18]<=1; R_b[22][19]<=0;   
             R_b[23][0]<=0; R_b[23][1]<=0; R_b[23][2]<=0; R_b[23][3]<=0; R_b[23][4]<=1; R_b[23][5]<=1; R_b[23][6]<=0; R_b[23][7]<=0; R_b[23][8]<=0; R_b[23][9]<=0;R_b[23][10]<=0; R_b[23][11]<=0; R_b[23][12]<=1; R_b[23][13]<=1; R_b[23][14]<=1; R_b[23][15]<=1; R_b[23][16]<=1; R_b[23][17]<=0; R_b[23][18]<=0; R_b[23][19]<=0;
             R_b[24][0]<=0; R_b[24][1]<=0; R_b[24][2]<=0; R_b[24][3]<=0; R_b[24][4]<=0; R_b[24][5]<=0; R_b[24][6]<=0; R_b[24][7]<=0; R_b[24][8]<=0; R_b[24][9]<=1;R_b[24][10]<=1; R_b[24][11]<=0; R_b[24][12]<=1; R_b[24][13]<=0; R_b[24][14]<=0; R_b[24][15]<=0; R_b[24][16]<=1; R_b[24][17]<=0; R_b[24][18]<=0; R_b[24][19]<=0;
             R_b[25][0]<=1; R_b[25][1]<=1; R_b[25][2]<=1; R_b[25][3]<=0; R_b[25][4]<=0; R_b[25][5]<=0; R_b[25][6]<=0; R_b[25][7]<=0; R_b[25][8]<=0; R_b[25][9]<=0;R_b[25][10]<=0; R_b[25][11]<=0; R_b[25][12]<=1; R_b[25][13]<=0; R_b[25][14]<=0; R_b[25][15]<=0; R_b[25][16]<=1; R_b[25][17]<=0; R_b[25][18]<=0; R_b[25][19]<=0;
             R_b[26][0]<=0; R_b[26][1]<=0; R_b[26][2]<=1; R_b[26][3]<=0; R_b[26][4]<=0; R_b[26][5]<=0; R_b[26][6]<=0; R_b[26][7]<=0; R_b[26][8]<=0; R_b[26][9]<=0;R_b[26][10]<=0; R_b[26][11]<=0; R_b[26][12]<=1; R_b[26][13]<=0; R_b[26][14]<=0; R_b[26][15]<=0; R_b[26][16]<=1; R_b[26][17]<=0; R_b[26][18]<=0; R_b[26][19]<=0;
             R_b[27][0]<=0; R_b[27][1]<=0; R_b[27][2]<=1; R_b[27][3]<=1; R_b[27][4]<=1; R_b[27][5]<=1; R_b[27][6]<=0; R_b[27][7]<=1; R_b[27][8]<=0; R_b[27][9]<=0;R_b[27][10]<=0; R_b[27][11]<=0; R_b[27][12]<=0; R_b[27][13]<=0; R_b[27][14]<=0; R_b[27][15]<=0; R_b[27][16]<=1; R_b[27][17]<=0; R_b[27][18]<=0; R_b[27][19]<=0;
             R_b[28][0]<=0; R_b[28][1]<=0; R_b[28][2]<=0; R_b[28][3]<=0; R_b[28][4]<=0; R_b[28][5]<=1; R_b[28][6]<=0; R_b[28][7]<=0; R_b[28][8]<=1; R_b[28][9]<=0;R_b[28][10]<=0; R_b[28][11]<=0; R_b[28][12]<=0; R_b[28][13]<=0; R_b[28][14]<=0; R_b[28][15]<=0; R_b[28][16]<=0; R_b[28][17]<=0; R_b[28][18]<=0; R_b[28][19]<=0;
             R_b[29][0]<=0; R_b[29][1]<=0; R_b[29][2]<=0; R_b[29][3]<=0; R_b[29][4]<=0; R_b[29][5]<=1; R_b[29][6]<=0; R_b[29][7]<=0; R_b[29][8]<=0; R_b[29][9]<=1;R_b[29][10]<=1; R_b[29][11]<=1; R_b[29][12]<=1; R_b[29][13]<=1; R_b[29][14]<=0; R_b[29][15]<=0; R_b[29][16]<=0; R_b[29][17]<=0; R_b[29][18]<=1; R_b[29][19]<=0;
             R_b[30][0]<=0; R_b[30][1]<=0; R_b[30][2]<=0; R_b[30][3]<=0; R_b[30][4]<=0; R_b[30][5]<=0; R_b[30][6]<=0; R_b[30][7]<=0; R_b[30][8]<=0; R_b[30][9]<=0;R_b[30][10]<=0; R_b[30][11]<=0; R_b[30][12]<=0; R_b[30][13]<=0; R_b[30][14]<=0; R_b[30][15]<=0; R_b[30][16]<=0; R_b[30][17]<=0; R_b[30][18]<=1; R_b[30][19]<=0;   
             R_b[31][0]<=1; R_b[31][1]<=1; R_b[31][2]<=0; R_b[31][3]<=0; R_b[31][4]<=0; R_b[31][5]<=0; R_b[31][6]<=0; R_b[31][7]<=1; R_b[31][8]<=1; R_b[31][9]<=0;R_b[31][10]<=0; R_b[31][11]<=0; R_b[31][12]<=0; R_b[31][13]<=0; R_b[31][14]<=1; R_b[31][15]<=1; R_b[31][16]<=0; R_b[31][17]<=0; R_b[31][18]<=1; R_b[31][19]<=0;
             R_b[32][0]<=0; R_b[32][1]<=0; R_b[32][2]<=0; R_b[32][3]<=0; R_b[32][4]<=0; R_b[32][5]<=0; R_b[32][6]<=0; R_b[32][7]<=0; R_b[32][8]<=0; R_b[32][9]<=0;R_b[32][10]<=0; R_b[32][11]<=0; R_b[32][12]<=0; R_b[32][13]<=0; R_b[32][14]<=0; R_b[32][15]<=0; R_b[32][16]<=0; R_b[32][17]<=0; R_b[32][18]<=1; R_b[32][19]<=0;   
             R_b[33][0]<=0; R_b[33][1]<=0; R_b[33][2]<=0; R_b[33][3]<=0; R_b[33][4]<=1; R_b[33][5]<=1; R_b[33][6]<=1; R_b[33][7]<=0; R_b[33][8]<=0; R_b[33][9]<=0;R_b[33][10]<=1; R_b[33][11]<=1; R_b[33][12]<=1; R_b[33][13]<=1; R_b[33][14]<=1; R_b[33][15]<=0; R_b[33][16]<=0; R_b[33][17]<=0; R_b[33][18]<=1; R_b[33][19]<=0;
             R_b[34][0]<=0; R_b[34][1]<=0; R_b[34][2]<=0; R_b[34][3]<=0; R_b[34][4]<=0; R_b[34][5]<=0; R_b[34][6]<=0; R_b[34][7]<=0; R_b[34][8]<=0; R_b[34][9]<=0;R_b[34][10]<=0; R_b[34][11]<=0; R_b[34][12]<=0; R_b[34][13]<=0; R_b[34][14]<=0; R_b[34][15]<=0; R_b[34][16]<=0; R_b[34][17]<=0; R_b[34][18]<=1; R_b[34][19]<=0;
             R_b[35][0]<=0; R_b[35][1]<=0; R_b[35][2]<=1; R_b[35][3]<=0; R_b[35][4]<=0; R_b[35][5]<=0; R_b[35][6]<=0; R_b[35][7]<=1; R_b[35][8]<=0; R_b[35][9]<=0;R_b[35][10]<=0; R_b[35][11]<=0; R_b[35][12]<=0; R_b[35][13]<=0; R_b[35][14]<=0; R_b[35][15]<=1; R_b[35][16]<=1; R_b[35][17]<=1; R_b[35][18]<=1; R_b[35][19]<=0;
             R_b[36][0]<=0; R_b[36][1]<=0; R_b[36][2]<=0; R_b[36][3]<=1; R_b[36][4]<=0; R_b[36][5]<=0; R_b[36][6]<=1; R_b[36][7]<=0; R_b[36][8]<=0; R_b[36][9]<=0;R_b[36][10]<=0; R_b[36][11]<=0; R_b[36][12]<=0; R_b[36][13]<=0; R_b[36][14]<=0; R_b[36][15]<=0; R_b[36][16]<=0; R_b[36][17]<=0; R_b[36][18]<=0; R_b[36][19]<=0;
             R_b[37][0]<=0; R_b[37][1]<=0; R_b[37][2]<=0; R_b[37][3]<=0; R_b[37][4]<=1; R_b[37][5]<=1; R_b[37][6]<=0; R_b[37][7]<=0; R_b[37][8]<=0; R_b[37][9]<=1;R_b[37][10]<=0; R_b[37][11]<=0; R_b[37][12]<=1; R_b[37][13]<=0; R_b[37][14]<=0; R_b[37][15]<=0; R_b[37][16]<=0; R_b[37][17]<=0; R_b[37][18]<=0; R_b[37][19]<=0;
             R_b[38][0]<=1; R_b[38][1]<=1; R_b[38][2]<=0; R_b[38][3]<=0; R_b[38][4]<=0; R_b[38][5]<=0; R_b[38][6]<=0; R_b[38][7]<=0; R_b[38][8]<=0; R_b[38][9]<=1;R_b[38][10]<=0; R_b[38][11]<=0; R_b[38][12]<=1; R_b[38][13]<=0; R_b[38][14]<=0; R_b[38][15]<=0; R_b[38][16]<=0; R_b[38][17]<=0; R_b[38][18]<=0; R_b[38][19]<=1;
             R_b[39][0]<=0; R_b[39][1]<=0; R_b[39][2]<=0; R_b[39][3]<=0; R_b[39][4]<=0; R_b[39][5]<=0; R_b[39][6]<=0; R_b[39][7]<=0; R_b[39][8]<=0; R_b[39][9]<=0;R_b[39][10]<=0; R_b[39][11]<=0; R_b[39][12]<=1; R_b[39][13]<=1; R_b[39][14]<=1; R_b[39][15]<=1; R_b[39][16]<=1; R_b[39][17]<=0; R_b[39][18]<=0; R_b[39][19]<=1;             
            end                
        else if (store)
        begin
             R_b[n][m]<=1;
             //R_b[n_r1][m_r1]<=0;
             R_b[n_r2][m_r2]<=0;
            // R_b[n_r3][m_r3]<=0;
             //R_b[n_r4][m_r4]<=0;
        end
      end
    
 always @ (posedge clk or posedge clr)
    begin   
        if (clr)
            begin 
            //01 /1 19/  8 15/ 24 13/  29 8 / 35 6
             R_q[0][0]<=0; R_q[0][1]<=1; R_q[0][2]<=0; R_q[0][3]<=0; R_q[0][4]<=0; R_q[0][5]<=0; R_q[0][6]<=0; R_q[0][7]<=0; R_q[0][8]<=0; R_q[0][9]<=0;R_q[0][10]<=0; R_q[0][11]<=0; R_q[0][12]<=0; R_q[0][13]<=0; R_q[0][14]<=0; R_q[0][15]<=0; R_q[0][16]<=0; R_q[0][17]<=0; R_q[0][18]<=0; R_q[0][19]<=0;
             R_q[1][0]<=0; R_q[1][1]<=0; R_q[1][2]<=0; R_q[1][3]<=0; R_q[1][4]<=0; R_q[1][5]<=0; R_q[1][6]<=0; R_q[1][7]<=0; R_q[1][8]<=0; R_q[1][9]<=0;R_q[1][10]<=0; R_q[1][11]<=0; R_q[1][12]<=0; R_q[1][13]<=0; R_q[1][14]<=0; R_q[1][15]<=0; R_q[1][16]<=0; R_q[1][17]<=0; R_q[1][18]<=0; R_q[1][19]<=0;
             R_q[2][0]<=0; R_q[2][1]<=0; R_q[2][2]<=0; R_q[2][3]<=0; R_q[2][4]<=0; R_q[2][5]<=0; R_q[2][6]<=0; R_q[2][7]<=0; R_q[2][8]<=0; R_q[2][9]<=0;R_q[2][10]<=0; R_q[2][11]<=0; R_q[2][12]<=0; R_q[2][13]<=0; R_q[2][14]<=0; R_q[2][15]<=0; R_q[2][16]<=0; R_q[2][17]<=0; R_q[2][18]<=0; R_q[2][19]<=0;
             R_q[3][0]<=0; R_q[3][1]<=0; R_q[3][2]<=0; R_q[3][3]<=0; R_q[3][4]<=0; R_q[3][5]<=0; R_q[3][6]<=0; R_q[3][7]<=0; R_q[3][8]<=0; R_q[3][9]<=0;R_q[3][10]<=0; R_q[3][11]<=0; R_q[3][12]<=0; R_q[3][13]<=0; R_q[3][14]<=0; R_q[3][15]<=0; R_q[3][16]<=0; R_q[3][17]<=0; R_q[3][18]<=0; R_q[3][19]<=0;
             R_q[4][0]<=0; R_q[4][1]<=0; R_q[4][2]<=0; R_q[4][3]<=0; R_q[4][4]<=0; R_q[4][5]<=0; R_q[4][6]<=0; R_q[4][7]<=0; R_q[4][8]<=0; R_q[4][9]<=0;R_q[4][10]<=0; R_q[4][11]<=0; R_q[4][12]<=0; R_q[4][13]<=0; R_q[4][14]<=0; R_q[4][15]<=0; R_q[4][16]<=0; R_q[4][17]<=0; R_q[4][18]<=0; R_q[4][19]<=0;
             R_q[5][0]<=0; R_q[5][1]<=0; R_q[5][2]<=0; R_q[5][3]<=0; R_q[5][4]<=0; R_q[5][5]<=0; R_q[5][6]<=0; R_q[5][7]<=0; R_q[5][8]<=0; R_q[5][9]<=0;R_q[5][10]<=0; R_q[5][11]<=0; R_q[5][12]<=0; R_q[5][13]<=0; R_q[5][14]<=0; R_q[5][15]<=0; R_q[5][16]<=0; R_q[5][17]<=0; R_q[5][18]<=0; R_q[5][19]<=0;
             R_q[6][0]<=0; R_q[6][1]<=0; R_q[6][2]<=0; R_q[6][3]<=0; R_q[6][4]<=0; R_q[6][5]<=0; R_q[6][6]<=0; R_q[6][7]<=0; R_q[6][8]<=0; R_q[6][9]<=0;R_q[6][10]<=0; R_q[6][11]<=0; R_q[6][12]<=0; R_q[6][13]<=0; R_q[6][14]<=0; R_q[6][15]<=0; R_q[6][16]<=0; R_q[6][17]<=0; R_q[6][18]<=0; R_q[6][19]<=0;           
             R_q[7][0]<=0; R_q[7][1]<=0; R_q[7][2]<=0; R_q[7][3]<=0; R_q[7][4]<=0; R_q[7][5]<=0; R_q[7][6]<=0; R_q[7][7]<=0; R_q[7][8]<=0; R_q[7][9]<=0;R_q[7][10]<=0; R_q[7][11]<=0; R_q[7][12]<=0; R_q[7][13]<=0; R_q[7][14]<=0; R_q[7][15]<=0; R_q[7][16]<=0; R_q[7][17]<=0; R_q[7][18]<=0; R_q[7][19]<=0;   
             R_q[8][0]<=0; R_q[8][1]<=0; R_q[8][2]<=0; R_q[8][3]<=0; R_q[8][4]<=0; R_q[8][5]<=0; R_q[8][6]<=0; R_q[8][7]<=0; R_q[8][8]<=0; R_q[8][9]<=0;R_q[8][10]<=0; R_q[8][11]<=0; R_q[8][12]<=0; R_q[8][13]<=0; R_q[8][14]<=0; R_q[8][15]<=0; R_q[8][16]<=0; R_q[8][17]<=0; R_q[8][18]<=0; R_q[8][19]<=0;   
             R_q[9][0]<=0; R_q[9][1]<=0; R_q[9][2]<=0; R_q[9][3]<=0; R_q[9][4]<=0; R_q[9][5]<=0; R_q[9][6]<=0; R_q[9][7]<=0; R_q[9][8]<=0; R_q[9][9]<=0;R_q[9][10]<=0; R_q[9][11]<=0; R_q[9][12]<=0; R_q[9][13]<=0; R_q[9][14]<=0; R_q[9][15]<=0; R_q[9][16]<=0; R_q[9][17]<=0; R_q[9][18]<=0; R_q[9][19]<=0;   
             R_q[10][0]<=0; R_q[10][1]<=0; R_q[10][2]<=0; R_q[10][3]<=0; R_q[10][4]<=0; R_q[10][5]<=0; R_q[10][6]<=0; R_q[10][7]<=0; R_q[10][8]<=0; R_q[10][9]<=0;R_q[10][10]<=0; R_q[10][11]<=0; R_q[10][12]<=0; R_q[10][13]<=0; R_q[10][14]<=0; R_q[10][15]<=0; R_q[10][16]<=0; R_q[10][17]<=0; R_q[10][18]<=0; R_q[10][19]<=0;   
             R_q[11][0]<=0; R_q[11][1]<=0; R_q[11][2]<=0; R_q[11][3]<=0; R_q[11][4]<=0; R_q[11][5]<=0; R_q[11][6]<=0; R_q[11][7]<=0; R_q[11][8]<=0; R_q[11][9]<=0;R_q[11][10]<=0; R_q[11][11]<=0; R_q[11][12]<=0; R_q[11][13]<=0; R_q[11][14]<=0; R_q[11][15]<=0; R_q[11][16]<=0; R_q[11][17]<=0; R_q[11][18]<=0; R_q[11][19]<=0;
             R_q[12][0]<=0; R_q[12][1]<=0; R_q[12][2]<=0; R_q[12][3]<=0; R_q[12][4]<=0; R_q[12][5]<=0; R_q[12][6]<=0; R_q[12][7]<=0; R_q[12][8]<=0; R_q[12][9]<=0;R_q[12][10]<=0; R_q[12][11]<=0; R_q[12][12]<=0; R_q[12][13]<=0; R_q[12][14]<=0; R_q[12][15]<=0; R_q[12][16]<=0; R_q[12][17]<=0; R_q[12][18]<=0; R_q[12][19]<=0;   
             R_q[13][0]<=0; R_q[13][1]<=0; R_q[13][2]<=0; R_q[13][3]<=0; R_q[13][4]<=0; R_q[13][5]<=0; R_q[13][6]<=0; R_q[13][7]<=0; R_q[13][8]<=0; R_q[13][9]<=0;R_q[13][10]<=0; R_q[13][11]<=0; R_q[13][12]<=0; R_q[13][13]<=0; R_q[13][14]<=0; R_q[13][15]<=0; R_q[13][16]<=0; R_q[13][17]<=0; R_q[13][18]<=0; R_q[13][19]<=0;
             R_q[14][0]<=0; R_q[14][1]<=0; R_q[14][2]<=0; R_q[14][3]<=0; R_q[14][4]<=0; R_q[14][5]<=0; R_q[14][6]<=0; R_q[14][7]<=0; R_q[14][8]<=0; R_q[14][9]<=0;R_q[14][10]<=0; R_q[14][11]<=0; R_q[14][12]<=0; R_q[14][13]<=0; R_q[14][14]<=0; R_q[14][15]<=0; R_q[14][16]<=0; R_q[14][17]<=0; R_q[14][18]<=0; R_q[14][19]<=0;
             R_q[15][0]<=0; R_q[15][1]<=0; R_q[15][2]<=0; R_q[15][3]<=0; R_q[15][4]<=0; R_q[15][5]<=0; R_q[15][6]<=0; R_q[15][7]<=0; R_q[15][8]<=0; R_q[15][9]<=0;R_q[15][10]<=0; R_q[15][11]<=0; R_q[15][12]<=0; R_q[15][13]<=0; R_q[15][14]<=0; R_q[15][15]<=0; R_q[15][16]<=0; R_q[15][17]<=0; R_q[15][18]<=0; R_q[15][19]<=0;
             R_q[16][0]<=0; R_q[16][1]<=0; R_q[16][2]<=0; R_q[16][3]<=0; R_q[16][4]<=0; R_q[16][5]<=0; R_q[16][6]<=0; R_q[16][7]<=0; R_q[16][8]<=0; R_q[16][9]<=0;R_q[16][10]<=0; R_q[16][11]<=0; R_q[16][12]<=0; R_q[16][13]<=0; R_q[16][14]<=0; R_q[16][15]<=0; R_q[16][16]<=0; R_q[16][17]<=0; R_q[16][18]<=0; R_q[16][19]<=0;
             R_q[17][0]<=0; R_q[17][1]<=0; R_q[17][2]<=0; R_q[17][3]<=0; R_q[17][4]<=0; R_q[17][5]<=0; R_q[17][6]<=0; R_q[17][7]<=0; R_q[17][8]<=0; R_q[17][9]<=0;R_q[17][10]<=0; R_q[17][11]<=0; R_q[17][12]<=0; R_q[17][13]<=0; R_q[17][14]<=0; R_q[17][15]<=0; R_q[17][16]<=0; R_q[17][17]<=0; R_q[17][18]<=0; R_q[17][19]<=0;
             R_q[18][0]<=0; R_q[18][1]<=0; R_q[18][2]<=0; R_q[18][3]<=0; R_q[18][4]<=0; R_q[18][5]<=0; R_q[18][6]<=0; R_q[18][7]<=0; R_q[18][8]<=0; R_q[18][9]<=0;R_q[18][10]<=0; R_q[18][11]<=0; R_q[18][12]<=0; R_q[18][13]<=0; R_q[18][14]<=0; R_q[18][15]<=0; R_q[18][16]<=0; R_q[18][17]<=0; R_q[18][18]<=0; R_q[18][19]<=0;
             R_q[19][0]<=0; R_q[19][1]<=0; R_q[19][2]<=0; R_q[19][3]<=0; R_q[19][4]<=0; R_q[19][5]<=0; R_q[19][6]<=0; R_q[19][7]<=0; R_q[19][8]<=0; R_q[19][9]<=0;R_q[19][10]<=0; R_q[19][11]<=0; R_q[19][12]<=0; R_q[19][13]<=0; R_q[19][14]<=0; R_q[19][15]<=0; R_q[19][16]<=0; R_q[19][17]<=0; R_q[19][18]<=0; R_q[19][19]<=0;
             R_q[20][0]<=0; R_q[20][1]<=0; R_q[20][2]<=0; R_q[20][3]<=0; R_q[20][4]<=0; R_q[20][5]<=0; R_q[20][6]<=0; R_q[20][7]<=0; R_q[20][8]<=0; R_q[20][9]<=0;R_q[20][10]<=0; R_q[20][11]<=0; R_q[20][12]<=0; R_q[20][13]<=0; R_q[20][14]<=0; R_q[20][15]<=0; R_q[20][16]<=0; R_q[20][17]<=0; R_q[20][18]<=0; R_q[20][19]<=0;   
             R_q[21][0]<=0; R_q[21][1]<=0; R_q[21][2]<=0; R_q[21][3]<=0; R_q[21][4]<=0; R_q[21][5]<=0; R_q[21][6]<=0; R_q[21][7]<=0; R_q[21][8]<=0; R_q[21][9]<=0;R_q[21][10]<=0; R_q[21][11]<=0; R_q[21][12]<=0; R_q[21][13]<=0; R_q[21][14]<=0; R_q[21][15]<=0; R_q[21][16]<=0; R_q[21][17]<=0; R_q[21][18]<=0; R_q[21][19]<=0;
             R_q[22][0]<=0; R_q[22][1]<=0; R_q[22][2]<=0; R_q[22][3]<=0; R_q[22][4]<=0; R_q[22][5]<=0; R_q[22][6]<=0; R_q[22][7]<=0; R_q[22][8]<=0; R_q[22][9]<=0;R_q[22][10]<=0; R_q[22][11]<=0; R_q[22][12]<=0; R_q[22][13]<=0; R_q[22][14]<=0; R_q[22][15]<=0; R_q[22][16]<=0; R_q[22][17]<=0; R_q[22][18]<=0; R_q[22][19]<=0;   
             R_q[23][0]<=0; R_q[23][1]<=0; R_q[23][2]<=0; R_q[23][3]<=0; R_q[23][4]<=0; R_q[23][5]<=0; R_q[23][6]<=0; R_q[23][7]<=0; R_q[23][8]<=0; R_q[23][9]<=0;R_q[23][10]<=0; R_q[23][11]<=0; R_q[23][12]<=0; R_q[23][13]<=0; R_q[23][14]<=0; R_q[23][15]<=0; R_q[23][16]<=0; R_q[23][17]<=0; R_q[23][18]<=0; R_q[23][19]<=0;
             R_q[24][0]<=0; R_q[24][1]<=0; R_q[24][2]<=0; R_q[24][3]<=0; R_q[24][4]<=0; R_q[24][5]<=0; R_q[24][6]<=0; R_q[24][7]<=0; R_q[24][8]<=0; R_q[24][9]<=0;R_q[24][10]<=0; R_q[24][11]<=0; R_q[24][12]<=0; R_q[24][13]<=0; R_q[24][14]<=0; R_q[24][15]<=0; R_q[24][16]<=0; R_q[24][17]<=0; R_q[24][18]<=0; R_q[24][19]<=0;
             R_q[25][0]<=0; R_q[25][1]<=0; R_q[25][2]<=0; R_q[25][3]<=0; R_q[25][4]<=0; R_q[25][5]<=0; R_q[25][6]<=0; R_q[25][7]<=0; R_q[25][8]<=0; R_q[25][9]<=0;R_q[25][10]<=0; R_q[25][11]<=0; R_q[25][12]<=0; R_q[25][13]<=0; R_q[25][14]<=0; R_q[25][15]<=0; R_q[25][16]<=0; R_q[25][17]<=0; R_q[25][18]<=0; R_q[25][19]<=0;
             R_q[26][0]<=0; R_q[26][1]<=0; R_q[26][2]<=0; R_q[26][3]<=0; R_q[26][4]<=0; R_q[26][5]<=0; R_q[26][6]<=0; R_q[26][7]<=0; R_q[26][8]<=0; R_q[26][9]<=0;R_q[26][10]<=0; R_q[26][11]<=0; R_q[26][12]<=0; R_q[26][13]<=0; R_q[26][14]<=0; R_q[26][15]<=0; R_q[26][16]<=0; R_q[26][17]<=0; R_q[26][18]<=0; R_q[26][19]<=0;
             R_q[27][0]<=0; R_q[27][1]<=0; R_q[27][2]<=0; R_q[27][3]<=0; R_q[27][4]<=0; R_q[27][5]<=0; R_q[27][6]<=0; R_q[27][7]<=0; R_q[27][8]<=0; R_q[27][9]<=0;R_q[27][10]<=0; R_q[27][11]<=0; R_q[27][12]<=0; R_q[27][13]<=0; R_q[27][14]<=0; R_q[27][15]<=0; R_q[27][16]<=0; R_q[27][17]<=0; R_q[27][18]<=0; R_q[27][19]<=0;
             R_q[28][0]<=0; R_q[28][1]<=0; R_q[28][2]<=0; R_q[28][3]<=0; R_q[28][4]<=0; R_q[28][5]<=0; R_q[28][6]<=0; R_q[28][7]<=0; R_q[28][8]<=0; R_q[28][9]<=0;R_q[28][10]<=0; R_q[28][11]<=0; R_q[28][12]<=0; R_q[28][13]<=0; R_q[28][14]<=0; R_q[28][15]<=0; R_q[28][16]<=0; R_q[28][17]<=0; R_q[28][18]<=0; R_q[28][19]<=0;
             R_q[29][0]<=0; R_q[29][1]<=0; R_q[29][2]<=0; R_q[29][3]<=0; R_q[29][4]<=0; R_q[29][5]<=0; R_q[29][6]<=0; R_q[29][7]<=0; R_q[29][8]<=0; R_q[29][9]<=0;R_q[29][10]<=0; R_q[29][11]<=0; R_q[29][12]<=0; R_q[29][13]<=0; R_q[29][14]<=0; R_q[29][15]<=0; R_q[29][16]<=0; R_q[29][17]<=0; R_q[29][18]<=0; R_q[29][19]<=0;
             R_q[30][0]<=0; R_q[30][1]<=0; R_q[30][2]<=0; R_q[30][3]<=0; R_q[30][4]<=0; R_q[30][5]<=0; R_q[30][6]<=0; R_q[30][7]<=0; R_q[30][8]<=0; R_q[30][9]<=0;R_q[30][10]<=0; R_q[30][11]<=0; R_q[30][12]<=0; R_q[30][13]<=0; R_q[30][14]<=0; R_q[30][15]<=0; R_q[30][16]<=0; R_q[30][17]<=0; R_q[30][18]<=0; R_q[30][19]<=0;   
             R_q[31][0]<=0; R_q[31][1]<=0; R_q[31][2]<=0; R_q[31][3]<=0; R_q[31][4]<=0; R_q[31][5]<=0; R_q[31][6]<=0; R_q[31][7]<=0; R_q[31][8]<=0; R_q[31][9]<=0;R_q[31][10]<=0; R_q[31][11]<=0; R_q[31][12]<=0; R_q[31][13]<=0; R_q[31][14]<=0; R_q[31][15]<=0; R_q[31][16]<=0; R_q[31][17]<=0; R_q[31][18]<=0; R_q[31][19]<=0;
             R_q[32][0]<=0; R_q[32][1]<=0; R_q[32][2]<=0; R_q[32][3]<=0; R_q[32][4]<=0; R_q[32][5]<=0; R_q[32][6]<=0; R_q[32][7]<=0; R_q[32][8]<=0; R_q[32][9]<=0;R_q[32][10]<=0; R_q[32][11]<=0; R_q[32][12]<=0; R_q[32][13]<=0; R_q[32][14]<=0; R_q[32][15]<=0; R_q[32][16]<=0; R_q[32][17]<=0; R_q[32][18]<=0; R_q[32][19]<=0;   
             R_q[33][0]<=0; R_q[33][1]<=0; R_q[33][2]<=0; R_q[33][3]<=0; R_q[33][4]<=0; R_q[33][5]<=0; R_q[33][6]<=0; R_q[33][7]<=0; R_q[33][8]<=0; R_q[33][9]<=0;R_q[33][10]<=0; R_q[33][11]<=0; R_q[33][12]<=0; R_q[33][13]<=0; R_q[33][14]<=0; R_q[33][15]<=0; R_q[33][16]<=0; R_q[33][17]<=0; R_q[33][18]<=0; R_q[33][19]<=0;
             R_q[34][0]<=0; R_q[34][1]<=0; R_q[34][2]<=0; R_q[34][3]<=0; R_q[34][4]<=0; R_q[34][5]<=0; R_q[34][6]<=0; R_q[34][7]<=0; R_q[34][8]<=0; R_q[34][9]<=0;R_q[34][10]<=0; R_q[34][11]<=0; R_q[34][12]<=0; R_q[34][13]<=0; R_q[34][14]<=0; R_q[34][15]<=0; R_q[34][16]<=0; R_q[34][17]<=0; R_q[34][18]<=0; R_q[34][19]<=0;
             R_q[35][0]<=0; R_q[35][1]<=0; R_q[35][2]<=0; R_q[35][3]<=0; R_q[35][4]<=0; R_q[35][5]<=0; R_q[35][6]<=0; R_q[35][7]<=0; R_q[35][8]<=0; R_q[35][9]<=0;R_q[35][10]<=0; R_q[35][11]<=0; R_q[35][12]<=0; R_q[35][13]<=0; R_q[35][14]<=0; R_q[35][15]<=0; R_q[35][16]<=0; R_q[35][17]<=0; R_q[35][18]<=0; R_q[35][19]<=0;
             R_q[36][0]<=0; R_q[36][1]<=0; R_q[36][2]<=0; R_q[36][3]<=0; R_q[36][4]<=0; R_q[36][5]<=0; R_q[36][6]<=0; R_q[36][7]<=0; R_q[36][8]<=0; R_q[36][9]<=0;R_q[36][10]<=0; R_q[36][11]<=0; R_q[36][12]<=0; R_q[36][13]<=0; R_q[36][14]<=0; R_q[36][15]<=0; R_q[36][16]<=0; R_q[36][17]<=0; R_q[36][18]<=0; R_q[36][19]<=0;
             R_q[37][0]<=0; R_q[37][1]<=0; R_q[37][2]<=0; R_q[37][3]<=0; R_q[37][4]<=0; R_q[37][5]<=0; R_q[37][6]<=0; R_q[37][7]<=0; R_q[37][8]<=0; R_q[37][9]<=0;R_q[37][10]<=0; R_q[37][11]<=0; R_q[37][12]<=0; R_q[37][13]<=0; R_q[37][14]<=0; R_q[37][15]<=0; R_q[37][16]<=0; R_q[37][17]<=0; R_q[37][18]<=0; R_q[37][19]<=0;
             R_q[38][0]<=0; R_q[38][1]<=0; R_q[38][2]<=0; R_q[38][3]<=0; R_q[38][4]<=0; R_q[38][5]<=0; R_q[38][6]<=0; R_q[38][7]<=0; R_q[38][8]<=0; R_q[38][9]<=0;R_q[38][10]<=0; R_q[38][11]<=0; R_q[38][12]<=0; R_q[38][13]<=0; R_q[38][14]<=0; R_q[38][15]<=0; R_q[38][16]<=0; R_q[38][17]<=0; R_q[38][18]<=0; R_q[38][19]<=0;
             R_q[39][0]<=0; R_q[39][1]<=0; R_q[39][2]<=0; R_q[39][3]<=0; R_q[39][4]<=0; R_q[39][5]<=0; R_q[39][6]<=0; R_q[39][7]<=0; R_q[39][8]<=0; R_q[39][9]<=0;R_q[39][10]<=0; R_q[39][11]<=0; R_q[39][12]<=0; R_q[39][13]<=0; R_q[39][14]<=0; R_q[39][15]<=0; R_q[39][16]<=0; R_q[39][17]<=0; R_q[39][18]<=0; R_q[39][19]<=0; 
           end
       else if (store)
        begin
             R_q[n][m]<=0;
             end
           end
           
 always@(*) 
    begin       
      if (judge)
        begin
            if ((|R_q[0])|(|R_q[1])|(|R_q[2])|(|R_q[3])|(|R_q[4])|(|R_q[5])|(|R_q[6])|(|R_q[7])|(|R_q[8])|(|R_q[9])|(|R_q[10])|(|R_q[11])|(|R_q[12])|(|R_q[13])|(|R_q[14])|(|R_q[15])|(|R_q[16])|(|R_q[17])|(|R_q[18])|(|R_q[19])|(|R_q[20])|(|R_q[21])|(|R_q[22])|(|R_q[23])|(|R_q[24])|(|R_q[25])|(|R_q[26])|(|R_q[27])|(|R_q[28])|(|R_q[29])|(|R_q[30])|(|R_q[31])|(|R_q[32])|(|R_q[33])|(|R_q[34])|(|R_q[35])|(|R_q[36])|(|R_q[37])|(|R_q[38])  |(|R_q[39]))
                judge_able=0;
            end
            else if(!((|R_q[0])|(|R_q[1])|(|R_q[2])|(|R_q[3])|(|R_q[4])|(|R_q[5])|(|R_q[6])|(|R_q[7])|(|R_q[8])|(|R_q[9])|(|R_q[10])|(|R_q[11])|(|R_q[12])|(|R_q[13])|(|R_q[14])|(|R_q[15])|(|R_q[16])|(|R_q[17])|(|R_q[18])|(|R_q[19])|(|R_q[20])|(|R_q[21])|(|R_q[22])|(|R_q[23])|(|R_q[24])|(|R_q[25])|(|R_q[26])|(|R_q[27])|(|R_q[28])|(|R_q[29])|(|R_q[30])|(|R_q[31])|(|R_q[32])|(|R_q[33])|(|R_q[34])|(|R_q[35])|(|R_q[36])|(|R_q[37])|(|R_q[38])  |(|R_q[39])))
                 judge_able=1;
    end

 
 always @ (posedge clk or posedge clr)
    begin
        if (clr)
            n <= 0;
        else if ((move_able==1)&&(d_r==1))
            n <= n+1;
        else if ((move_able==1)&&(u_r==1))
            n <= n-1;
        else
            n <= n;
    end
  
  always @ (posedge clk or posedge clr)
    begin
        if (clr)
            m <= 0;
        else if  ((move_able==1)&&(l_r==1))
             m <= m-1;
        else if  ((move_able==1)&&(r_r==1))
             m <= m+1;
        else
            m <= m;
    end
                          
endmodule
